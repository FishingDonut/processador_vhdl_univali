--by Daniel Uesler de Brito.
-- Trabalho em trios, mas todos devem saber explicar o projeto inteiro.

-- Consulte o guia prático do risc-v para entender sobre o formato das instruções.
---- conecte os campos das instruções no processador
------ exemplo: separando os 7 bits de opcode da instrução w_INST(6 downto 0)



-- Crie um módulo controle
---- A interface do controle está comentada neste documento.
---- Gere os sinais de controle de acordo com o código de operação recebido.
---- Ligue os sinais corretamente.
---- DICA: Saber como esses sinais funcionam garante uma questão da prova.



-- Modifique a ULA para receber o sinal de w_ALUOP do controle.
---- Ele serve, entre outras coisas, para evitar que a ULA tente fazer uma operação de SUBI incorretamente.
---- A ULA deve realizar, pelo menos, as operações de ADD/SUB, AND, OR, XOR


-- Inclua a memória de dados e seu caminho de dados.
---- Com esse arquivo será possível fazer operações de LW e SW.
---- A memória de dados deve receber: 
------ A saída w_ULA como entrada de endereço.
------ A saída w_RS2 como entrada de dados.
------ Controlar a operação com sinais do controle.

-- Inclua um multiplexador no projeto para que o controle possa escolher entre colocar o dado que sai da ULA ou da memória de dados no banco de registradores


-- Não é necessário implementar o caminho dos desvios condicionais e incondicionais, mas é desejável que o controle gere o sinal de desvio

-- OBS: 
---- Seu código só vai começar a compilar quando você conectar os sinais que estão em aberto no código.
---- Você terá que modificar a memória de instruções para testar operações de LW e SW
---- Utilizem o simulador da Cadence em Tools & Simulators, pois ele executa o diagrama de formas de onda corretamente.



library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity RISCV32i is

	Port (	i_CLK  	: in  std_logic;
    		i_RSTn	: in  std_logic;
            
            -- sinais de para depuração
            o_INST		: out std_logic_vector(31 downto 0);
            o_OPCODE	: out std_logic_vector(6 downto 0);
            o_RD_ADDR	: out std_logic_vector(4 downto 0);
            o_RS1_ADDR 	: out std_logic_vector(4 downto 0);
            o_RS2_ADDR 	: out std_logic_vector(4 downto 0);
            o_RS1_DATA 	: out std_logic_vector(31 downto 0);
            o_RS2_DATA 	: out std_logic_vector(31 downto 0);
            o_IMM   	: out std_logic_vector(31 downto 0);
            o_ULA   	: out std_logic_vector(31 downto 0);
            o_MEM   	: out std_logic_vector(31 downto 0)
         );

end RISCV32i;

architecture arch_1 of RISCV32i is
	signal w_RS1, w_RS2 : std_logic_vector(31 downto 0); -- liga a saída do banco
    signal w_ULA : std_logic_vector(31 downto 0); -- liga a saída da ULA
    signal w_ULAb: std_logic_vector(31 downto 0); -- liga entrada b da ula
    signal w_ZERO: std_logic; 
    
    --sinais da memória de dados
    signal w_MEM: std_logic_vector(31 downto 0); -- saída da memória de dados
    
    -- sinais do gerador de imediato
    signal w_IMM : std_logic_vector(31 downto 0);
    -- sinais do pc e memória de instrução
    signal w_PC, w_PC4 : std_logic_vector(31 downto 0); -- endereço da instrução/ próxima instrução
    signal w_INST : std_logic_vector(31 downto 0); -- instrução lida
    
    -- sinais de controle
    signal w_ALU_SRC	: std_logic;
    signal w_MEM2REG	: std_logic;
    signal w_REG_WRITE	: std_logic;
    signal w_MEM_READ	: std_logic;
    signal w_MEM_WRITE	: std_logic;
    signal w_ALUOP    	: std_logic_vector(1 downto 0);
    
begin

    
    

	u_CONTROLE: entity work.controle
	port map (	
    	i_OPCODE 	=> w_INST(6 downto 0),
    	o_ALU_SRC	=> w_ALU_SRC, -- escolhe entre w_RS2 e w_IMED
        o_MEM2REG	=> w_MEM2REG, -- escolhe entre w_ALU e w_MEM
        o_REG_WRITE	=> w_REG_WRITE, -- permite escrever no BANCO DE REGISTRADORES
        o_MEM_READ	=> w_MEM_READ, -- habilita memória para leitura
        o_MEM_WRITE	=> w_MEM_WRITE, -- habilita memória para escrita
        o_ALUOP    	=> w_ALUOP	-- gera sinais para ajudar a escolher a operação da ULA
    );

	u_PC: entity work.ffd -- registra o PC (próxima instrução a ser executada) 
    port map (
        i_DATA    => w_PC4, 
        i_CLK     => i_CLK,
        i_RSTn    => i_RSTn,
        o_DATA    => w_PC
    );
    
    u_SOMA4 : entity work.somador -- calcula o endereço da próxima instrução
	port map (	
    	i_A		=> w_PC, 
    	i_B  	=> "00000000000000000000000000000100",  
        o_DATA  => w_PC4
    );
    
	u_MEM_INST: entity work.memoria_instrucoes
    port map(
        i_ADDR		=> w_PC,
        o_INST 		=> w_INST
    );
    
    u_GERADOR_IMM : entity work.gerador_imediato -- gera o imediato concatenando os bits corretos (ext de sinal)
    port map(
        i_INST	=> w_INST,
        o_IMM   => w_IMM
    );

	u_BANCO_REGISTRADORES: entity work.banco_registradores
      port map (	
          i_CLK  	=> i_CLK, 
          i_RSTn	=> i_RSTn, 
          i_WRena	=> , -- coloque os campos corretos do controle
          i_WRaddr  => , -- coloque os campos corretos da instrução
          i_RS1 	=> , -- coloque os campos corretos da instrução
          i_RS2 	=> , -- coloque os campos corretos da instrução
          i_DATA 	=> w_ULA, 
          o_RS1 	=> w_RS1,	
          o_RS2 	=> w_RS2	
	);

	u_ULA : entity work.ULA 
    port map(
        i_A   	=> w_RS1,
        i_B   	=> w_ULAb,
        i_F3  	=> , -- coloque os campos corretos da instrução
        i_INST30=> , -- coloque os campos corretos da instrução
        o_ZERO   => w_ZERO, 
        o_ULA => w_ULA
    );
    
    u_MUX_ULA: entity work.mux21
    port map (
    	i_A		=> w_RS2, 
        i_B		=> , -- coloque os campos corretos da extensão de sinal
        i_SEL	=> , -- coloque os campos corretos do controle
        o_MUX   => w_ULAb 
    );
    
    --Sinais para depuração com o testbench
    o_INST 		<= w_INST; -- depuração do resultado da ula
    o_OPCODE	<= w_INST(6 downto 0);
    o_RD_ADDR	<= w_INST(11 downto 7);
    o_RS1_ADDR 	<= w_INST(19 downto 15);
    o_RS2_ADDR 	<= w_INST(24 downto 20);
    o_RS1_DATA 	<= w_RS1;
    o_RS2_DATA 	<= w_RS2;
    o_IMM   	<= w_IMM;
    o_ULA 		<= w_ULA; -- depuração do resultado da ula
    o_MEM		<= w_MEM;
    



end arch_1;